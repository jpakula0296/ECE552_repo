module cache_arbiter(
  input [15:0] instr_addr, instr_cache_in, data_addr, data_cache_in,
  input instr_miss, data_miss,

  output memory_address

);



endmodule
