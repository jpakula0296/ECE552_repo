module cpu(
  input clk, rst_n,
  output hlt,
  output [15:0] pc
  );
