module IF_ID(
    input [15:0] instr_in,
    input [15:0] pc_current_in
    output [15:0] instr_out,
    output [15:0] pc_current_out
    );
