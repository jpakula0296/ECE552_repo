module cache_block_decoder(
  input [6:0] block_num,
  output reg [127:0] BlockEnable
);

reg [127:0] BlockEnable;
wire [127:0] base;
assign base = 127'h1; // shift this left to get values

// implementing with shifts so we don't have to type out all these values
always @* case(shift_val)
7'd0 : BlockEnable = base << 7'd0;
7'd1 : BlockEnable = base << 7'd1;
7'd2 : BlockEnable = base << 7'd2;
7'd3 : BlockEnable = base << 7'd3;
7'd4 : BlockEnable = base << 7'd4;
7'd5 : BlockEnable = base << 7'd5;
7'd6 : BlockEnable = base << 7'd6;
7'd7 : BlockEnable = base << 7'd7;
7'd8 : BlockEnable = base << 7'd8;
7'd9 : BlockEnable = base << 7'd9;
7'd10 : BlockEnable = base << 7'd10;
7'd11 : BlockEnable = base << 7'd11;
7'd12 : BlockEnable = base << 7'd12;
7'd13 : BlockEnable = base << 7'd13;
7'd14 : BlockEnable = base << 7'd14;
7'd15 : BlockEnable = base << 7'd15;
7'd16 : BlockEnable = base << 7'd16;
7'd17 : BlockEnable = base << 7'd17;
7'd18 : BlockEnable = base << 7'd18;
7'd19 : BlockEnable = base << 7'd19;
7'd20 : BlockEnable = base << 7'd20;
7'd21 : BlockEnable = base << 7'd21;
7'd22 : BlockEnable = base << 7'd22;
7'd23 : BlockEnable = base << 7'd23;
7'd24 : BlockEnable = base << 7'd24;
7'd25 : BlockEnable = base << 7'd25;
7'd26 : BlockEnable = base << 7'd26;
7'd27 : BlockEnable = base << 7'd27;
7'd28 : BlockEnable = base << 7'd28;
7'd29 : BlockEnable = base << 7'd29;
7'd30 : BlockEnable = base << 7'd30;
7'd31 : BlockEnable = base << 7'd31;
7'd32 : BlockEnable = base << 7'd32;
7'd33 : BlockEnable = base << 7'd33;
7'd34 : BlockEnable = base << 7'd34;
7'd35 : BlockEnable = base << 7'd35;
7'd36 : BlockEnable = base << 7'd36;
7'd37 : BlockEnable = base << 7'd37;
7'd38 : BlockEnable = base << 7'd38;
7'd39 : BlockEnable = base << 7'd39;
7'd40 : BlockEnable = base << 7'd40;
7'd41 : BlockEnable = base << 7'd41;
7'd42 : BlockEnable = base << 7'd42;
7'd43 : BlockEnable = base << 7'd43;
7'd44 : BlockEnable = base << 7'd44;
7'd45 : BlockEnable = base << 7'd45;
7'd46 : BlockEnable = base << 7'd46;
7'd47 : BlockEnable = base << 7'd47;
7'd48 : BlockEnable = base << 7'd48;
7'd49 : BlockEnable = base << 7'd49;
7'd50 : BlockEnable = base << 7'd50;
7'd51 : BlockEnable = base << 7'd51;
7'd52 : BlockEnable = base << 7'd52;
7'd53 : BlockEnable = base << 7'd53;
7'd54 : BlockEnable = base << 7'd54;
7'd55 : BlockEnable = base << 7'd55;
7'd56 : BlockEnable = base << 7'd56;
7'd57 : BlockEnable = base << 7'd57;
7'd58 : BlockEnable = base << 7'd58;
7'd59 : BlockEnable = base << 7'd59;
7'd60 : BlockEnable = base << 7'd60;
7'd61 : BlockEnable = base << 7'd61;
7'd62 : BlockEnable = base << 7'd62;
7'd63 : BlockEnable = base << 7'd63;
7'd64 : BlockEnable = base << 7'd64;
7'd65 : BlockEnable = base << 7'd65;
7'd66 : BlockEnable = base << 7'd66;
7'd67 : BlockEnable = base << 7'd67;
7'd68 : BlockEnable = base << 7'd68;
7'd69 : BlockEnable = base << 7'd69;
7'd70 : BlockEnable = base << 7'd70;
7'd71 : BlockEnable = base << 7'd71;
7'd72 : BlockEnable = base << 7'd72;
7'd73 : BlockEnable = base << 7'd73;
7'd74 : BlockEnable = base << 7'd74;
7'd75 : BlockEnable = base << 7'd75;
7'd76 : BlockEnable = base << 7'd76;
7'd77 : BlockEnable = base << 7'd77;
7'd78 : BlockEnable = base << 7'd78;
7'd79 : BlockEnable = base << 7'd79;
7'd80 : BlockEnable = base << 7'd80;
7'd81 : BlockEnable = base << 7'd81;
7'd82 : BlockEnable = base << 7'd82;
7'd83 : BlockEnable = base << 7'd83;
7'd84 : BlockEnable = base << 7'd84;
7'd85 : BlockEnable = base << 7'd85;
7'd86 : BlockEnable = base << 7'd86;
7'd87 : BlockEnable = base << 7'd87;
7'd88 : BlockEnable = base << 7'd88;
7'd89 : BlockEnable = base << 7'd89;
7'd90 : BlockEnable = base << 7'd90;
7'd91 : BlockEnable = base << 7'd91;
7'd92 : BlockEnable = base << 7'd92;
7'd93 : BlockEnable = base << 7'd93;
7'd94 : BlockEnable = base << 7'd94;
7'd95 : BlockEnable = base << 7'd95;
7'd96 : BlockEnable = base << 7'd96;
7'd97 : BlockEnable = base << 7'd97;
7'd98 : BlockEnable = base << 7'd98;
7'd99 : BlockEnable = base << 7'd99;
7'd100 : BlockEnable = base << 7'd100;
7'd101 : BlockEnable = base << 7'd101;
7'd102 : BlockEnable = base << 7'd102;
7'd103 : BlockEnable = base << 7'd103;
7'd104 : BlockEnable = base << 7'd104;
7'd105 : BlockEnable = base << 7'd105;
7'd106 : BlockEnable = base << 7'd106;
7'd107 : BlockEnable = base << 7'd107;
7'd108 : BlockEnable = base << 7'd108;
7'd109 : BlockEnable = base << 7'd109;
7'd110 : BlockEnable = base << 7'd110;
7'd111 : BlockEnable = base << 7'd111;
7'd112 : BlockEnable = base << 7'd112;
7'd113 : BlockEnable = base << 7'd113;
7'd114 : BlockEnable = base << 7'd114;
7'd115 : BlockEnable = base << 7'd115;
7'd116 : BlockEnable = base << 7'd116;
7'd117 : BlockEnable = base << 7'd117;
7'd118 : BlockEnable = base << 7'd118;
7'd119 : BlockEnable = base << 7'd119;
7'd120 : BlockEnable = base << 7'd120;
7'd121 : BlockEnable = base << 7'd121;
7'd122 : BlockEnable = base << 7'd122;
7'd123 : BlockEnable = base << 7'd123;
7'd124 : BlockEnable = base << 7'd124;
7'd125 : BlockEnable = base << 7'd125;
7'd126 : BlockEnable = base << 7'd126;
7'd127 : BlockEnable = base << 7'd127;



endmodule
