module full_adder(
  input A,
  input B,
  input Cin,

  output Sum,
  output Cout;
  );
