module MEM_data(
    input [15:0] ALU_Out_in,
    input [15:0] rt_in,
    input data_wr_in,
    output [15:0] ALU_Out_out,
    output [15:0] rt_in,
    output data_wr_in,
);
endmodule
