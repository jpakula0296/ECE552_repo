module WriteDecoder_4_16(
  input [3:0] RegId,
  input WriteReg,
  output [15:0] Wordline
  );

  
