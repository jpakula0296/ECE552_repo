module 4bit_Ripple_Carry_tb();
