module addsub_4bit_tb();
