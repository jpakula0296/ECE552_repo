module BitCell(
  input clk, rst, D, WriteEnable, ReadEnable1, ReadEnable2,
  inout Bitline1, Bitline2
  );
  
