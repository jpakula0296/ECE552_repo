/*
 * 16 bit ALU, capable of performing the following operations:
 *      ADD
 *      PADDSB
 *      SUB
 *      XOR
 *      RED
 *      SLL
 *      SRA
 *      ROR
 */
module alu(
    input [15:0]    rs,
    input [15:0]    rt,
    output [15:0]   rd,
);
endmodule
