module MEM_data(
    input [15:0] ALU_Out,
    input [15:0] rt,
    input data_wr,
);
endmodule
