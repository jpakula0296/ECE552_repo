module ID_data(
    input [15:0] instr_in,
    input [15:0] pc_plus_four_in,
    output [15:0] instr_out,
    output [15:0] pc_plus_four_out
    );
