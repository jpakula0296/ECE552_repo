module addsub_4bit( );
