module cache_block_decoder(
  input [6:0] block_num,
  output [127:0] BlockEnable
);

reg [127:0] BlockEnable_reg;
wire [127:0] base;
assign base = 127'h1; // shift this left to get values
assign BlockEnable = BlockEnable_reg;

// implementing with shifts so we don't have to type out all these values
always @* case(block_num)
7'd0 : BlockEnable_reg = base << 7'd0;
7'd1 : BlockEnable_reg = base << 7'd1;
7'd2 : BlockEnable_reg = base << 7'd2;
7'd3 : BlockEnable_reg = base << 7'd3;
7'd4 : BlockEnable_reg = base << 7'd4;
7'd5 : BlockEnable_reg = base << 7'd5;
7'd6 : BlockEnable_reg = base << 7'd6;
7'd7 : BlockEnable_reg = base << 7'd7;
7'd8 : BlockEnable_reg = base << 7'd8;
7'd9 : BlockEnable_reg = base << 7'd9;
7'd10 : BlockEnable_reg = base << 7'd10;
7'd11 : BlockEnable_reg = base << 7'd11;
7'd12 : BlockEnable_reg = base << 7'd12;
7'd13 : BlockEnable_reg = base << 7'd13;
7'd14 : BlockEnable_reg = base << 7'd14;
7'd15 : BlockEnable_reg = base << 7'd15;
7'd16 : BlockEnable_reg = base << 7'd16;
7'd17 : BlockEnable_reg = base << 7'd17;
7'd18 : BlockEnable_reg = base << 7'd18;
7'd19 : BlockEnable_reg = base << 7'd19;
7'd20 : BlockEnable_reg = base << 7'd20;
7'd21 : BlockEnable_reg = base << 7'd21;
7'd22 : BlockEnable_reg = base << 7'd22;
7'd23 : BlockEnable_reg = base << 7'd23;
7'd24 : BlockEnable_reg = base << 7'd24;
7'd25 : BlockEnable_reg = base << 7'd25;
7'd26 : BlockEnable_reg = base << 7'd26;
7'd27 : BlockEnable_reg = base << 7'd27;
7'd28 : BlockEnable_reg = base << 7'd28;
7'd29 : BlockEnable_reg = base << 7'd29;
7'd30 : BlockEnable_reg = base << 7'd30;
7'd31 : BlockEnable_reg = base << 7'd31;
7'd32 : BlockEnable_reg = base << 7'd32;
7'd33 : BlockEnable_reg = base << 7'd33;
7'd34 : BlockEnable_reg = base << 7'd34;
7'd35 : BlockEnable_reg = base << 7'd35;
7'd36 : BlockEnable_reg = base << 7'd36;
7'd37 : BlockEnable_reg = base << 7'd37;
7'd38 : BlockEnable_reg = base << 7'd38;
7'd39 : BlockEnable_reg = base << 7'd39;
7'd40 : BlockEnable_reg = base << 7'd40;
7'd41 : BlockEnable_reg = base << 7'd41;
7'd42 : BlockEnable_reg = base << 7'd42;
7'd43 : BlockEnable_reg = base << 7'd43;
7'd44 : BlockEnable_reg = base << 7'd44;
7'd45 : BlockEnable_reg = base << 7'd45;
7'd46 : BlockEnable_reg = base << 7'd46;
7'd47 : BlockEnable_reg = base << 7'd47;
7'd48 : BlockEnable_reg = base << 7'd48;
7'd49 : BlockEnable_reg = base << 7'd49;
7'd50 : BlockEnable_reg = base << 7'd50;
7'd51 : BlockEnable_reg = base << 7'd51;
7'd52 : BlockEnable_reg = base << 7'd52;
7'd53 : BlockEnable_reg = base << 7'd53;
7'd54 : BlockEnable_reg = base << 7'd54;
7'd55 : BlockEnable_reg = base << 7'd55;
7'd56 : BlockEnable_reg = base << 7'd56;
7'd57 : BlockEnable_reg = base << 7'd57;
7'd58 : BlockEnable_reg = base << 7'd58;
7'd59 : BlockEnable_reg = base << 7'd59;
7'd60 : BlockEnable_reg = base << 7'd60;
7'd61 : BlockEnable_reg = base << 7'd61;
7'd62 : BlockEnable_reg = base << 7'd62;
7'd63 : BlockEnable_reg = base << 7'd63;
7'd64 : BlockEnable_reg = base << 7'd64;
7'd65 : BlockEnable_reg = base << 7'd65;
7'd66 : BlockEnable_reg = base << 7'd66;
7'd67 : BlockEnable_reg = base << 7'd67;
7'd68 : BlockEnable_reg = base << 7'd68;
7'd69 : BlockEnable_reg = base << 7'd69;
7'd70 : BlockEnable_reg = base << 7'd70;
7'd71 : BlockEnable_reg = base << 7'd71;
7'd72 : BlockEnable_reg = base << 7'd72;
7'd73 : BlockEnable_reg = base << 7'd73;
7'd74 : BlockEnable_reg = base << 7'd74;
7'd75 : BlockEnable_reg = base << 7'd75;
7'd76 : BlockEnable_reg = base << 7'd76;
7'd77 : BlockEnable_reg = base << 7'd77;
7'd78 : BlockEnable_reg = base << 7'd78;
7'd79 : BlockEnable_reg = base << 7'd79;
7'd80 : BlockEnable_reg = base << 7'd80;
7'd81 : BlockEnable_reg = base << 7'd81;
7'd82 : BlockEnable_reg = base << 7'd82;
7'd83 : BlockEnable_reg = base << 7'd83;
7'd84 : BlockEnable_reg = base << 7'd84;
7'd85 : BlockEnable_reg = base << 7'd85;
7'd86 : BlockEnable_reg = base << 7'd86;
7'd87 : BlockEnable_reg = base << 7'd87;
7'd88 : BlockEnable_reg = base << 7'd88;
7'd89 : BlockEnable_reg = base << 7'd89;
7'd90 : BlockEnable_reg = base << 7'd90;
7'd91 : BlockEnable_reg = base << 7'd91;
7'd92 : BlockEnable_reg = base << 7'd92;
7'd93 : BlockEnable_reg = base << 7'd93;
7'd94 : BlockEnable_reg = base << 7'd94;
7'd95 : BlockEnable_reg = base << 7'd95;
7'd96 : BlockEnable_reg = base << 7'd96;
7'd97 : BlockEnable_reg = base << 7'd97;
7'd98 : BlockEnable_reg = base << 7'd98;
7'd99 : BlockEnable_reg = base << 7'd99;
7'd100 : BlockEnable_reg = base << 7'd100;
7'd101 : BlockEnable_reg = base << 7'd101;
7'd102 : BlockEnable_reg = base << 7'd102;
7'd103 : BlockEnable_reg = base << 7'd103;
7'd104 : BlockEnable_reg = base << 7'd104;
7'd105 : BlockEnable_reg = base << 7'd105;
7'd106 : BlockEnable_reg = base << 7'd106;
7'd107 : BlockEnable_reg = base << 7'd107;
7'd108 : BlockEnable_reg = base << 7'd108;
7'd109 : BlockEnable_reg = base << 7'd109;
7'd110 : BlockEnable_reg = base << 7'd110;
7'd111 : BlockEnable_reg = base << 7'd111;
7'd112 : BlockEnable_reg = base << 7'd112;
7'd113 : BlockEnable_reg = base << 7'd113;
7'd114 : BlockEnable_reg = base << 7'd114;
7'd115 : BlockEnable_reg = base << 7'd115;
7'd116 : BlockEnable_reg = base << 7'd116;
7'd117 : BlockEnable_reg = base << 7'd117;
7'd118 : BlockEnable_reg = base << 7'd118;
7'd119 : BlockEnable_reg = base << 7'd119;
7'd120 : BlockEnable_reg = base << 7'd120;
7'd121 : BlockEnable_reg = base << 7'd121;
7'd122 : BlockEnable_reg = base << 7'd122;
7'd123 : BlockEnable_reg = base << 7'd123;
7'd124 : BlockEnable_reg = base << 7'd124;
7'd125 : BlockEnable_reg = base << 7'd125;
7'd126 : BlockEnable_reg = base << 7'd126;
7'd127 : BlockEnable_reg = base << 7'd127;
endcase

endmodule
