module PC_tb();

endmodule
